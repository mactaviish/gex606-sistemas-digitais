`include "pasta/mux.v"

module tarefa_5(entrada_x, resultado);
    reg [16:0] Reg_S, Reg_H;
    reg [8:0] Reg_X;
    mux m0, m1, m2;
    ula ula;

endmodule