module somador (input [3:0] a,b, output [3:0] res);
	assign res = a + b;
endmodule